* Pixel Circuit
.include p18_cmos_models_tt.inc
.include PhotoDiode.inc

.subckt PIXEL VDD VSS EXPOSE ERASE NRE OUT
	* Photodiode
	XPD1	N1	VDD	PhotoDiode
	
	* Expose trigger
	M1	N1 	EXPOSE 	N2	0 	NMOS 	L=LNswitch 	W=WNswitch
	
	* Erase trigger
	M2	N2	ERASE		0	0 	NMOS 	L=LNswitch 	W=WNswitch
	
	* Sampling Capacitor
	Cs	N2	0	3p
	
	* Readout circuit
	M3 	N3 	N2 	0 	VDD 	PMOS 	L=LPamp 	W=WPamp
	M4 	OUT 	NRE	N3 	VDD 	PMOS 	L=LPamp 	W=WPamp

.ends PIXEL