* Pixel Circuit
.include p18_cmos_models_tt.inc
.include PhotoDiode.inc

.subckt PIXEL VDD VSS EXPOSE ERASE NRE OUT
	* Parameters
	.param LN = 1U
	.param kN = 2
	.param WN = {kN*LN}
	
	.param LP = 1U
	.param kP = 7.14
	.param WP = {kP*LP}
	
	* Photodiode
	XPD1	VDD	N1	PhotoDiode
	
	* Expose trigger
	M1	N1 	EXPOSE 	N2	0 	NMOS 	L=LN 	W=WN
	
	* Erase trigger
	M2	N2	ERASE		0	0 	NMOS 	L=LN 	W=WN
	
	* Sampling Capacitor
	Cs	N2	0	10f
	
	* Readout circuit
	M3 	N3 	N2 	0 	VDD 	PMOS 	L=LP 	W=WP
	M4 	OUT 	NRE	N3 	VDD 	PMOS 	L=LP 	W=WP

.ends PIXEL