[aimspice]
[description]
1837
* Pixel testbench
.include pixel_circuit.cir

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

* Transistor Parameters ***********************
* NMOS Switches - tune for high closed impedance
.param LNswitch = 2U
.param WNswitch = 2U

* NMOS Switches - tune for low open impedance
.param LPswitch = 0.7U
.param WPswitch = 10U

* Amplifiers - tune for linearity
.param LPamp = 0.7U
.param WPamp = 10U

* Active loads - tune for linearity
.param LPload = 2U
.param WPload = 2U

**********************************

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE NRE 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)

* Photodiode
XPD1	1	N1	PhotoDiode	Ipd=550
	
* Expose trigger
M1	N1 	EXPOSE 	N2	0 	NMOS 	L=LNswitch 	W=WNswitch
	
* Erase trigger
M2	N2	ERASE		0	0	NMOS 	L=LNswitch 	W=WNswitch
	
* Sampling Capacitor
Cs	N2	0	3p
	
* Readout circuit
M3 	0 	N2 	N3 	1 	PMOS 	L=LPamp 	W=WPamp
M4 	N3 	NRE	OUT 	1 	PMOS 	L=LPswitch 	W=WPswitch
MC1 	OUT	OUT	1	1 	PMOS 	L=LPload	W=WPload
CC1	OUT	0	3p

VCS N2 0 dc 0

.plot V(OUT)
[options]
1
Gmin 1.0E-39
[dc]
1
VCS
0
1.8
0.05
[tran]
0.1ms
60ms
X
X
0
[ana]
1 0
[end]
