* Pixel array
.include pixel_circuit.cir

.subckt PIXELARRAY VDD VSS EXPOSE ERASE NRE_R1 NRE_R2 OUT1 OUT2
	* Pixels
	XP1_1 	VDD 	VSS 	EXPOSE 	ERASE 	NRE_R1 	OUT1	PIXEL
	XP1_2 	VDD 	VSS 	EXPOSE 	ERASE 	NRE_R1 	OUT2	PIXEL
	XP2_1 	VDD 	VSS 	EXPOSE 	ERASE 	NRE_R2 	OUT1	PIXEL
	XP2_2 	VDD 	VSS 	EXPOSE 	ERASE 	NRE_R2 	OUT2	PIXEL
	
	* Active loads 
	* Transistors
	MC1 	VDD	OUT1	OUT1	VDD 	PMOS 	L=LPload	W=WPload
	MC2 	VDD	OUT2	OUT2	VDD 	PMOS 	L=LPload	W=WPload
	* Parasitic Capacitors
	CC1	OUT1	0	3p
	CC2	OUT2	0	3p
	
.ends PIXELARRAY