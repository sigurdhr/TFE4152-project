[aimspice]
[description]
1455
* Pixel testbench
.include pixel_circuit.cir

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

* Transistor Parameters ***********************
.param LNswitch = 1U
.param kNswitch = 6
.param WNswitch = {kNswitch*LNswitch}
	
.param LPswitch = 1U
.param kPswitch = 6
.param WPswitch = {kPswitch*LPswitch}

.param LPamp = 1U
.param kPamp = 6
.param WPamp = {kPamp*LPamp}

.param LPload = 1U
.param kPload = 6
.param WPload = {kPload*LPload}

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VOUT OUT1 0 dc

XP1_1	1	0	EXPOSE	ERASE	NRE_R1	OUT1	PIXEL

.plot V(OUT1)
.plot V(EXPOSE) V(NRE_R1) V(ERASE)
[options]
1
Gmin 1.0E-39
[tran]
0.1ms
60ms
X
X
0
[ana]
4 0
[end]
