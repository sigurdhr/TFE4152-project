* Pixel array
.include pixel_circuit.cir

.subckt PIXELARRAY VDD VSSS EXPOSE ERASE NRE_R1 NRE_R2 OUT1 OUT2
	* Pixels
	XP1_1 	VDD 	VSSS 	EXPOSE 	ERASE 	NRE_R1 	OUT1	PIXEL	Ipd=Ipd_1
	XP1_2 	VDD 	VSSS 	EXPOSE 	ERASE 	NRE_R1 	OUT2	PIXEL	Ipd=Ipd_2	
	XP2_1 	VDD 	VSSS 	EXPOSE 	ERASE 	NRE_R2 	OUT1	PIXEL	Ipd=Ipd_3
	XP2_2 	VDD 	VSSS 	EXPOSE 	ERASE 	NRE_R2 	OUT2	PIXEL	Ipd=Ipd_4
	
	* Active loads 
	* Transistors
	MC1 	OUT1	OUT1	VDD	VDD 	PMOS 	L=LPload	W=WPload
	MC2 	OUT2	OUT2	VDD	VDD 	PMOS 	L=LPload	W=WPload
	* Parasitic Capacitors
	CC1	OUT1	0	3p
	CC2	OUT2	0	3p
	
.ends PIXELARRAY